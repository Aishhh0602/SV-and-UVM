interface fa_interface;
  logic a;
  logic b;
  logic cin;
  logic s;
  logic c;
  
endinterface